
hii from khaled