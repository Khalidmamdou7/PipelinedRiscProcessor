LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY CONTROL IS
PORT(
	clk : IN std_logic;
	OPcode : IN  std_logic_vector(4 DOWNTO 0);

	RegWrite : OUT std_logic;
    IOread : OUT std_logic;
    IOwrite : OUT std_logic;

    ISbranch : OUT std_logic;
    branchSRC : OUT std_logic_vector (1 DOWNTO 0);

    ALUoperation : OUT  std_logic_vector(2 DOWNTO 0);
    ALUSRC : OUT std_logic;

    Push : out std_logic;
    Pop : out std_logic;
    MemRead : out std_logic;
    MemWrite : out std_logic;

    RTI : out std_logic;
    RET : out std_logic;
    PCsrc2 : out std_logic;

    MemIndex : out std_logic_vector(1 DOWNTO 0);
    UseMemIndex : out std_logic;

    MemtoReg : out std_logic;

    selectorforCALL : out std_logic;
    selectorforINT : out std_logic
);
END ENTITY;

ARCHITECTURE myCONTROL OF CONTROL IS
	BEGIN
	PROCESS(clk) IS
		BEGIN
			if OPcode = "00000" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "11";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "00010" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "101";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "00011" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "010";
                ALUSRC <= '1';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "00100" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "011";
                ALUSRC <= '1';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "00101" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '1';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "00110" then
                RegWrite <= '0';
                IOread <= '1';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "00111" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "110";
                ALUSRC <= '1';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "01000" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "111";
                ALUSRC <= '1';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "01001" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "000";
                ALUSRC <= '1';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "01010" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "001";
                ALUSRC <= '1';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "01011" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "100";
                ALUSRC <= '1';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "01100" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "000";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "01110" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '1';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "01111" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '1';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "10000" then
                RegWrite <= '1';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "000";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '1';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "10001" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "00";
                ALUoperation <= "000";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '1';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "10010" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '1';
                branchSRC <= "00";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "10011" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '1';
                branchSRC <= "01";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "10100" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '1';
                branchSRC <= "10";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "10101" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '1';
                branchSRC <= "11";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '1';
                selectorforINT <= '1';
            elsif OPcode = "10110" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '1';
                branchSRC <= "11";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '1';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '0';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '0';
                selectorforINT <= '1';
            elsif OPcode = "10111" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "11";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '1';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '1';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '0';
                selectorforINT <= '0';
            elsif OPcode = "11000" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "11";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '1';
                Pop <= '0';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '0';
                RET <= '1';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '0';
                selectorforINT <= '0';
            elsif OPcode = "11001" then
                RegWrite <= '0';
                IOread <= '0';
                IOwrite <= '0';
                ISbranch <= '0';
                branchSRC <= "11";
                ALUoperation <= "110";
                ALUSRC <= '0';
                Push <= '0';
                Pop <= '1';
                MemRead <= '0';
                MemWrite <= '0';
                RTI <= '1';
                RET <= '1';
                PCsrc2 <= '0';
                MemIndex <= "00";
                UseMemIndex <= '0';
                MemtoReg <= '0';
                selectorforCALL <= '0';
                selectorforINT <= '0';
            end if;
	END PROCESS;
END Architecture;